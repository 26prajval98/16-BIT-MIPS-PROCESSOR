module instr_mem   
 (  
      input [15:0] pc,  
      output wire [15:0] instruction  
 );
      wire [3 : 0] rom_addr = pc[4 : 1];  
      reg [15:0] rom[15:0];  
      initial  
      begin  
                rom[0] = 16'b1110010010000000; //addi $1,$1,0  
                rom[1] = 16'b1110100100001010; //addi $2,$2,10
                rom[2] = 16'b1110110110000000; //addi $3,$3,0
                rom[3] = 16'b1111001000000001; //Loop:addi $4,$4,1
                rom[4] = 16'b1100100110000101; //beq $2,$3,exit
                rom[5] = 16'b0000010100010000; //add $1,$1,$2 
                rom[6] = 16'b0000101000100001; //sub $2,$2,$4  
                rom[7] = 16'b0100000000000100; //j loop 
                rom[8] = 16'b0000000000000000;  
                rom[9] = 16'b0000000000000000; 
                rom[10] = 16'b1111001000000111;//exit: addi $4,$4,7    
                rom[11] = 16'b0000000000000000;  
                rom[12] = 16'b0000000000000000;  
                rom[13] = 16'b0000000000000000;  
                rom[14] = 16'b0000000000000000;  
                rom[15] = 16'b0000000000000000;  
      end  
      assign instruction = (pc[15:0] < 32 )? rom[rom_addr[3:0]]: 16'd0;  
 endmodule 
